* SPICE3 file created from inv2.ext - technology: min2

.option scale=0.1u
* User needs to add below 2 lines*
.include NMOS-180nm.lib
.include PMOS-180nm.lib

M1000 out in vdd vdd pfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1001 out in gnd gnd nfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
C0 vdd out 0.18fF
C1 vdd in 0.07fF
C2 out gnd 0.05fF
C3 in gnd 0.19fF
C4 vdd gnd 0.41fF

* User needs to add below 2 lines*
Vdd vdd gnd 1.8
Vin in gnd pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10e-12 2e-09 0e-00
.control
run
.endc
.end

