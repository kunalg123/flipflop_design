magic
tech min2
timestamp 1559498764
<< nwell >>
rect -1 0 25 26
<< ntransistor >>
rect 11 -14 13 -6
<< ptransistor >>
rect 11 6 13 14
<< ndiffusion >>
rect 10 -14 11 -6
rect 13 -14 14 -6
<< pdiffusion >>
rect 10 6 11 14
rect 13 6 14 14
<< ndcontact >>
rect 6 -14 10 -6
rect 14 -14 18 -6
<< pdcontact >>
rect 6 6 10 14
rect 14 6 18 14
<< psubstratepcontact >>
rect 2 -23 6 -19
rect 10 -23 14 -19
rect 18 -23 22 -19
<< nsubstratencontact >>
rect 2 19 6 23
rect 10 19 14 23
rect 18 19 22 23
<< polysilicon >>
rect 11 14 13 17
rect 11 -2 13 6
rect 3 -4 13 -2
rect 11 -6 13 -4
rect 11 -17 13 -14
<< polycontact >>
rect -1 -5 3 -1
<< metal1 >>
rect 0 19 2 23
rect 6 14 10 23
rect 14 19 18 23
rect 22 19 24 23
rect 14 -1 18 6
rect -3 -5 -1 -1
rect 14 -5 22 -1
rect 14 -6 18 -5
rect 6 -23 10 -14
rect 14 -23 18 -19
<< labels >>
rlabel metal1 -3 -5 -3 -1 3 in
rlabel metal1 22 -5 22 -1 7 out
rlabel metal1 15 -22 15 -22 1 gnd!
rlabel metal1 23 20 23 20 7 vdd!
<< end >>
