magic
tech min2
timestamp 1559478838
<< nwell >>
rect -4 8 30 34
<< ntransistor >>
rect 8 -6 10 2
rect 16 -6 18 2
<< ptransistor >>
rect 8 14 10 22
rect 16 14 18 22
<< ndiffusion >>
rect 2 -2 3 2
rect 7 -2 8 2
rect 2 -6 8 -2
rect 10 -6 16 2
rect 18 -2 24 2
rect 18 -6 19 -2
rect 23 -6 24 -2
<< pdiffusion >>
rect 2 18 3 22
rect 7 18 8 22
rect 2 14 8 18
rect 10 18 16 22
rect 10 14 11 18
rect 15 14 16 18
rect 18 18 19 22
rect 23 18 24 22
rect 18 14 24 18
<< ndcontact >>
rect 3 -2 7 2
rect 19 -6 23 -2
<< pdcontact >>
rect 3 18 7 22
rect 11 14 15 18
rect 19 18 23 22
<< psubstratepcontact >>
rect 3 -15 7 -11
rect 11 -15 15 -11
rect 19 -15 23 -11
<< nsubstratencontact >>
rect 3 27 7 31
rect 11 27 15 31
rect 19 27 23 31
<< polysilicon >>
rect 8 22 10 25
rect 16 22 18 25
rect 8 2 10 14
rect 16 2 18 14
rect 8 -9 10 -6
rect 16 -9 18 -6
<< metal1 >>
rect 2 27 3 31
rect 7 27 11 31
rect 15 27 19 31
rect 23 27 24 31
rect 3 22 7 27
rect 19 22 23 27
rect 11 7 15 14
rect 3 4 15 7
rect 3 2 7 4
rect 19 -11 23 -6
rect 2 -15 3 -11
rect 7 -15 11 -11
rect 15 -15 19 -11
rect 23 -15 24 -11
<< labels >>
rlabel polysilicon 9 3 9 3 1 a
rlabel polysilicon 17 3 17 3 1 b
rlabel metal1 12 6 12 6 1 out
rlabel metal1 18 29 18 29 5 vdd!
rlabel metal1 17 -13 17 -13 1 gnd!
<< end >>
