* SPICE3 file created from nand1.ext - technology: min2

.option scale=0.1u
* User needs to add below 2 lines to include spice model files*
.include NMOS-180nm.lib
.include PMOS-180nm.lib

M1000 out a vdd vdd pfet w=8 l=2
+  ad=48 pd=28 as=96 ps=56
M1001 vdd b out vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_10_n6# a out gnd nfet w=8 l=2
+  ad=48 pd=28 as=48 ps=28
M1003 gnd b a_10_n6# gnd nfet w=8 l=2
+  ad=48 pd=28 as=0 ps=0
C0 vdd a 0.07fF
C1 vdd b 0.07fF
C2 vdd out 0.02fF
C3 a b 0.07fF
C4 a out 0.01fF
C5 out gnd 0.04fF
C6 b gnd 0.07fF
C7 a gnd 0.07fF
C8 vdd gnd 0.67fF


* User needs to add below lines for simulation*
Vdd vdd gnd 1.8
Va a gnd pulse(0 1.8 1p 10p 10p 1n 2n)
Vb b gnd pulse(0 1.8 1p 10p 10p 1.5n 3n)
.tran 10e-12 10e-09 0e-00
.control
run
.endc
.end


